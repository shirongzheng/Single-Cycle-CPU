LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BQE IS
	PORT(		SIGNAL SEL		: IN STD_LOGIC;
				QA_IN				: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				QB_IN				: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				PC					: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				SHIFT_2			: INOUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				EQUAL				: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
				INSTR				: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END BQE;

ARCHITECTURE STRUCTURE OF BQE IS
BEGIN
	PROCESS(SEL)
	BEGIN 
		IF(SEL = '1') THEN 
			EQUAL <= (NOT(QB_IN(15 DOWNTO 0) XOR QA_IN(15 DOWNTO 0)));
			IF(EQUAL = "1111111111111111") THEN
				SHIFT_2 <= TO_STDLOGICVECTOR(TO_BITVECTOR(QB_IN) SLL 2);
				INSTR <= STD_LOGIC_VECTOR(SIGNED(PC) + SIGNED(SHIFT_2(15 DOWNTO 0))+4);
			ELSIF	(EQUAL = "0000000000000000") THEN
				INSTR <= STD_LOGIC_VECTOR(UNSIGNED(PC)+4);
		ELSE INSTR <= STD_LOGIC_VECTOR(UNSIGNED(PC)+4);
			END IF;
		END IF;
	END PROCESS;
END STRUCTURE;