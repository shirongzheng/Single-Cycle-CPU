LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY OP_CONTROL_EXT IS
	PORT(		INSTR				: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				TO_ALU			: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
				IMMEDIATE_OUT	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				R_FORMAT			: OUT STD_LOGIC);
END OP_CONTROL_EXT;

ARCHITECTURE STRUCTURE OF OP_CONTROL_EXT IS
	SIGNAL OP			: STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL RS			: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL RT			: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL RD			: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL SHAMT	   : STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL FUNCT		: STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL IMMEDIATE	: STD_LOGIC_VECTOR(15 DOWNTO 0);
	
	BEGIN 
		PROCESS(INSTR)
		BEGIN 
			OP <= INSTR(31 DOWNTO 26);
			RS <= INSTR(25 DOWNTO 21);
			RT <= INSTR(20 DOWNTO 16);
			RD <= INSTR(15 DOWNTO 11);
			SHAMT <= INSTR(10 DOWNTO 6);
			FUNCT <= INSTR(5 DOWNTO 0);
			IMMEDIATE <= INSTR(15 DOWNTO 0);
			
			IF(OP = "000000") THEN TO_ALU <= "00";  --ADDITION
										  R_FORMAT <= '1';
				ELSIF (OP = "000001") THEN TO_ALU <= "01"; -- SUBTRACTION 
													R_FORMAT <= '1';
				ELSIF (OP = "000010") THEN TO_ALU <= "10"; --ORI
													R_FORMAT <= '0';
				IMMEDIATE_OUT <= X"0000" & IMMEDIATE;
			END IF;
		END PROCESS;
END STRUCTURE;