LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY direct_controller IS
	PORT(		DIR_ADDR 			: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				INSTRUCTION_REG	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				CONTROLLER			: IN STD_LOGIC:='0';
				OUT_ADDR				: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END direct_controller;

ARCHITECTURE Structure OF direct_controller IS
BEGIN 
	PROCESS(CONTROLLER) --Controller's process
		BEGIN
			IF (CONTROLLER = '1') THEN OUT_ADDR <= DIR_ADDR(4 DOWNTO 0);
				ELSE OUT_ADDR <= INSTRUCTION_REG(4 DOWNTO 0);
			END IF;
	END PROCESS;
END Structure;
