LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY WRITE_TO IS
	PORT(		
				OP 						: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				SIGNAL POWER			: IN STD_LOGIC;
				SIGNAL DIN				: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				SIGNAL PC_IN			: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				SIGNAL AIN				: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				SIGNAL DOUT				: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				SIGNAL PC				: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				SIGNAL ADDR_A			: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
				SIGNAL ADDR_B			: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
				SIGNAL WRITE_TO_ADDR	: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END WRITE_TO;

ARCHITECTURE STRUCTURE OF WRITE_TO IS 
BEGIN 
	PROCESS(POWER)
		BEGIN
			IF (POWER = '1') THEN
				CASE OP IS
					WHEN "0000" => DOUT(31 DOWNTO 28) <= DIN;
					WHEN "0001" => DOUT(27 DOWNTO 24) <= DIN;
					WHEN "0010" => DOUT(23 DOWNTO 20) <= DIN;
					WHEN "0011" => DOUT(19 DOWNTO 16) <= DIN;
					WHEN "0100" => DOUT(15 DOWNTO 12) <= DIN;
					WHEN "0101" => DOUT(11 DOWNTO 8) <= DIN;
					WHEN "0110" => DOUT(7 DOWNTO 4) <= DIN;
					WHEN "0111" => DOUT(3 DOWNTO 0) <= DIN;
					WHEN "1000" => ADDR_A <= AIN;
					WHEN "1001" => ADDR_B <= AIN;
					WHEN "1010" => WRITE_TO_ADDR <= AIN;
					WHEN "1110" => PC <= "00000000000000000000000000000000";
					WHEN "1111" => PC <= PC_IN;
					WHEN OTHERS => NULL;
				END CASE;
			END IF;
	END PROCESS;
END STRUCTURE;
				
					
					