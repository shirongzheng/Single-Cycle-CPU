LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RD_WR_32 IS
	PORT(		WR_RD				: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
				DIN				: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
				IN_ADDR			: IN STD_LOGIC_VECTOR(4  DOWNTO 0);
				DATA				: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				INSTRUCTIONS	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				OUT_ADDR			: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END RD_WR_32;

ARCHITECTURE Structure OF RD_WR_32 IS
BEGIN
		PROCESS(WR_RD)
			BEGIN 
				IF (WR_RD = "00") THEN DATA <= DIN(31 DOWNTO 0);
				ELSIF (WR_RD = "01") THEN OUT_ADDR <= IN_ADDR(4 DOWNTO 0);
				ELSIF (WR_RD = "10") THEN INSTRUCTIONS <= DIN(31 DOWNTO 0);
				END IF;
		END PROCESS;
END Structure;
		