LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ZERO_EXT IS 
	PORT(		SIGNAL OUTPUT		: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
				SIGNAL EXT16_32	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END ZERO_EXT;

ARCHITECTURE STRUCTURE OF ZERO_EXT IS
BEGIN 
	EXT16_32 <= "0000000000000000" & OUTPUT;
END STRUCTURE;